module timer
// Parameters section
#(
    parameter CLOCK_FREQ = 32'd5 // 50MHz frequency
)
// Ports section
(
    input        clk,
    input        rst_n,
    output [5:0] o_seconds,  // 0-59 seconds
    output [5:0] o_minutes,  // 0-59 minutes
    output [4:0] o_hours,     // 0-99 hours 
    output inc_day
);

  localparam ONE_SECOND = CLOCK_FREQ-1 ;  // (0-59 there are 60 clocks)

  // Internal logic 
  reg [ 5:0] seconds_cnt;  // 0-59 seconds
  reg [ 5:0] minutes_cnt;  // 0-59 minutes
  reg [ 6:0] hours_cnt;  // 0-99 hours (8'd99 is the maximum value possible on two 7seg digits)
  reg [31:0] counter_1sec;  // counts every clock cycle (max val is 2**32 > 4.2bln)
  reg inc_day_cnt;
  // Create the code for the Timer
  always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
      counter_1sec <= 0;
      seconds_cnt  <= 0;
      minutes_cnt  <= 0;
      hours_cnt    <= 0;
      inc_day_cnt  <=0;
    end else begin
      if (counter_1sec == ONE_SECOND) begin
        counter_1sec <= 0;

        if (seconds_cnt == 6'd59) begin  // increment the seconds counter
          seconds_cnt <= 0;

          if (minutes_cnt == 6'd59) begin  // increment the minutes counter
            minutes_cnt <= 0;

            if (hours_cnt == 5'd23) begin    // increment the hours counter (will roll over after 99 hours)						
              hours_cnt <= 0;
              inc_day_cnt  <=1;
            end else begin
              hours_cnt <= hours_cnt + 1'b1;
            end

          end else begin
            minutes_cnt <= minutes_cnt + 1'b1;
          end

        end else begin
          seconds_cnt <= seconds_cnt + 1'b1;
        end

      end else begin
        counter_1sec <= counter_1sec + 1'b1;
      end
    end
  end

  assign o_seconds = seconds_cnt;
  assign o_minutes = minutes_cnt;
  assign o_hours   = hours_cnt;
  assign inc_day   = inc_day_cnt;
endmodule

